`timescale 1ns / 1ps

module InstructionMemory(
    input [31:0] Address,                             // Input Address 
    output reg [31:0] Instruction); 

    reg [31:0] memory [0:1024];
    integer i;
    
    /* Please fill in the implementation here */
    initial begin 
    $readmemh("instructions.mem", memory);
    
    //$readmemh("instructions.mem",memory);
//      memory[0] <= 32'b00100000000010000000000000000000;	//	loop:	addi	$t0, $zero, 0
//memory[1] <= 32'b00000000000000000000000000000000;	//		nop
//memory[2] <= 32'b00000000000000000000000000000000;	//		nop
//memory[3] <= 32'b00000000000000000000000000000000;	//		nop
//memory[4] <= 32'b00000000000000000000000000000000;	//		nop
//memory[5] <= 32'b00000000000000000000000000000000;	//		nop
//memory[6] <= 32'b00100000000010010000000000000110;	//		addi	$t1, $zero, 6
//memory[7] <= 32'b00000000000000000000000000000000;	//		nop
//memory[8] <= 32'b00000000000000000000000000000000;	//		nop
//memory[9] <= 32'b00000000000000000000000000000000;	//		nop
//memory[10] <= 32'b00000000000000000000000000000000;	//		nop
//memory[11] <= 32'b00000000000000000000000000000000;	//		nop
//memory[12] <= 32'b00100000000010100000000000001010;	//		addi	$t2, $zero, 10
//memory[13] <= 32'b00000000000000000000000000000000;	//		nop
//memory[14] <= 32'b00000000000000000000000000000000;	//		nop
//memory[15] <= 32'b00000000000000000000000000000000;	//		nop
//memory[16] <= 32'b00000000000000000000000000000000;	//		nop
//memory[17] <= 32'b00000000000000000000000000000000;	//		nop
//memory[18] <= 32'b10101101000010010000000000000000;	//		sw	$t1, 0($t0)
//memory[19] <= 32'b00000000000000000000000000000000;	//		nop
//memory[20] <= 32'b00000000000000000000000000000000;	//		nop
//memory[21] <= 32'b00000000000000000000000000000000;	//		nop
//memory[22] <= 32'b00000000000000000000000000000000;	//		nop
//memory[23] <= 32'b00000000000000000000000000000000;	//		nop
//memory[24] <= 32'b10101101000010100000000000000100;	//		sw	$t2, 4($t0)
//memory[25] <= 32'b00000000000000000000000000000000;	//		nop
//memory[26] <= 32'b00000000000000000000000000000000;	//		nop
//memory[27] <= 32'b00000000000000000000000000000000;	//		nop
//memory[28] <= 32'b00000000000000000000000000000000;	//		nop
//memory[29] <= 32'b00000000000000000000000000000000;	//		nop
//memory[30] <= 32'b10001101000100000000000000000000;	//		lw	$s0, 0($t0)
//memory[31] <= 32'b00000000000000000000000000000000;	//		nop
//memory[32] <= 32'b00000000000000000000000000000000;	//		nop
//memory[33] <= 32'b00000000000000000000000000000000;	//		nop
//memory[34] <= 32'b00000000000000000000000000000000;	//		nop
//memory[35] <= 32'b00000000000000000000000000000000;	//		nop
//memory[36] <= 32'b10001101000100010000000000000100;	//		lw	$s1, 4($t0)
//memory[37] <= 32'b00000000000000000000000000000000;	//		nop
//memory[38] <= 32'b00000000000000000000000000000000;	//		nop
//memory[39] <= 32'b00000000000000000000000000000000;	//		nop
//memory[40] <= 32'b00000000000000000000000000000000;	//		nop
//memory[41] <= 32'b00000000000000000000000000000000;	//		nop
//memory[42] <= 32'b00000010001100000101100000100010;	//		sub	$t3, $s1, $s0
//memory[43] <= 32'b00000000000000000000000000000000;	//		nop
//memory[44] <= 32'b00000000000000000000000000000000;	//		nop
//memory[45] <= 32'b00000000000000000000000000000000;	//		nop
//memory[46] <= 32'b00000000000000000000000000000000;	//		nop
//memory[47] <= 32'b00000000000000000000000000000000;	//		nop
//memory[48] <= 32'b00000000000010110110000011000000;	//		sll	$t4, $t3, 3
//memory[49] <= 32'b00000000000000000000000000000000;	//		nop
//memory[50] <= 32'b00000000000000000000000000000000;	//		nop
//memory[51] <= 32'b00000000000000000000000000000000;	//		nop
//memory[52] <= 32'b00000000000000000000000000000000;	//		nop
//memory[53] <= 32'b00000000000000000000000000000000;	//		nop
//memory[54] <= 32'b00000000000011000110100010000010;	//		srl	$t5, $t4, 2
//memory[55] <= 32'b00000000000000000000000000000000;	//		nop
//memory[56] <= 32'b00000000000000000000000000000000;	//		nop
//memory[57] <= 32'b00000000000000000000000000000000;	//		nop
//memory[58] <= 32'b00000000000000000000000000000000;	//		nop
//memory[59] <= 32'b00000000000000000000000000000000;	//		nop
//memory[60] <= 32'b00001000000000000000000000000000;	//		j	loop
    end
    
//    assign Instruction = memory[Address>>2];
    
    always @ (Address) begin
        if (Address[0] == 0 && Address[1] == 0) begin
            Instruction <= memory[Address>>2];
        end
    end

endmodule